module NOT(
	input wire a,
	output wire c
);

assign c = ~a;

endmodule
